package pkg5 is
  constant c_invert : boolean;
end package pkg5;
