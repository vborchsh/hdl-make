module repro (input ia);
   wire       a;
   wire [0:31] s;

/*
  mygate inst (a);
 */
endmodule
