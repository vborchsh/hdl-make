module mygate(input d);
endmodule
