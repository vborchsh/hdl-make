entity gate4 is
  port (i : in bit;
        o : out bit);
end gate4;
