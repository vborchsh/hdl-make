architecture behav of gate4 is
begin
  inst: entity work.gate
    port map (i, o);
end behav;
