package body pkg5 is
  constant c_invert : boolean := true;
end package body pkg5;
